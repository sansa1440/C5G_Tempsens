//=======================================================
//	LCD Module
//	
//	Using material
//	SC2004CSWB-XA-LB-G	
//	VDD=3.3 V

//Source
//http://www.cs.hiroshima-u.ac.jp/~nakano/wiki/wiki.cgi?page=lcdctrl%2Ev
//=======================================================

`define INIT    2'b00
`define SETPOS0 2'b01
`define SETPOS1 2'b10 
`define WRITE   2'b11

module lcdctrl_init(
	clk,
	reset,
	lcd_e,
	lcd_rs,
	lcd_rw,
	sf_d,
	);
	
	input clk,reset;
	output lcd_e,lcd_rs,lcd_rw;
	output [11:8] sf_d;

	reg lcd_e;
	reg [1:0] state = `INIT;
	reg [2:0] index;
	reg [3:0] addr;
	reg [31:0] counter;
	reg [30:0] ctrl;
	reg [7:0] ascii;
	reg [3:0] hex;

	wire set_enb;
	wire ret;
	wire [19:0] wait_cnt;


	assign lcd_rw   = 0;
	assign ret      = ctrl[30];
	assign lcd_rs   = ctrl[29];
	assign set_enb  = ctrl[28];
	assign sf_d     = ctrl[27:20];
	assign wait_cnt = ctrl[19:0];

	
	always @(posedge clk or negedge reset)
		if(!reset) begin
			addr <= 0;
			counter <= 0;
			state <= `INIT;
			index <= 0;
		end else if(counter<wait_cnt)
			counter <= counter + 1;
		else begin
			counter <= 0;
			if(!ret)
				addr <= addr + 1;
			else begin
					addr <= 0;
				if(state==`INIT)
					state <= `SETPOS0;
				else if(state==`SETPOS0 || state==`SETPOS1)
					state <= `WRITE;
				else if(state == `WRITE) begin
					if(index== 5)
						index <= 0;
					else
						index <= index + 1;
					if(index == 2)
						state <= `SETPOS1;
					else if(index == 5)
						state <= `SETPOS0;
			end
		end
	end

	always @(posedge clk or negedge reset) begin
		if(!reset) lcd_e <= 0;
		else if(set_enb && counter >= 1 && counter <= 12) lcd_e <= 1;
		else lcd_e <= 0;
	end

	always @(state or addr or ascii) begin
	case(state)
		`INIT:
		case(addr)
				4'h0: ctrl = {3'b000, 8'h00, 20'h03500};
				4'h1: ctrl = {3'b001, 8'h30, 20'h00550};
				4'h2: ctrl = {3'b001, 8'h30, 20'h00550};
				4'h3: ctrl = {3'b001, 8'h80, 20'h00550};
				4'h4: ctrl = {3'b101, 4'h00, 20'hF0800};
			default: ctrl = {3'bxxx, 8'h0x, 20'hxxxxx};
		endcase
//	`SETPOS0:
//	case(addr)
//	4'h0: ctrl = {3'b001, 4'h8, 20'h00041};
//	4'h1: ctrl = {3'b101, 4'h0, 20'h00800};
//	default: ctrl = {3'bxxx, 4'hx, 20'hxxxxx};
//	endcase
//	`SETPOS1:
//	case(addr)
//	4'h0 : ctrl = {3'b001, 4'hC, 20'h00041};
//	4'h1 : ctrl = {3'b101, 4'h0, 20'h00800};
//	default: ctrl = {3'bxxx, 4'hx, 20'hxxxxx};
//	endcase
//	`WRITE:
//	case(addr)
//	4'h0 : ctrl = {3'b011, ascii[7:4], 20'h00041};
//	4'h1 : ctrl = {3'b011, ascii[3:0], 20'h00800};
//	4'h2 : ctrl = {3'b011, ascii[7:4], 20'h00041};
//	4'h3 : ctrl = {3'b011, ascii[3:0], 20'h00800};
//	4'h4 : ctrl = {3'b011, ascii[7:4], 20'h00041};
//	4'h5 : ctrl = {3'b011, ascii[3:0], 20'h00800};
//	4'h6 : ctrl = {3'b011, ascii[7:4], 20'h00041};
//	4'h7 : ctrl = {3'b011, ascii[3:0], 20'h00800};
//	4'h8 : ctrl = {3'b011, 4'hA, 20'h00041};
//	4'h9 : ctrl = {3'b111, 4'h0, 20'h00800};
//	default: ctrl = {3'bxxx, 4'hx, 20'hxxxxx};
//	endcase
//	default: ctrl = {3'bxxx, 4'hx, 20'hxxxxx};
	endcase
	end

endmodule